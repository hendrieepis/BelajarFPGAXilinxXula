--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   20:24:14 02/26/2013
-- Design Name:   
-- Module Name:   /home/hendri/Documents/workspaceXilinx/keyboard_ps2/keybtest1.vhd
-- Project Name:  keyboard_ps2
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: keyboard
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;

entity keybtest1 is
end keybtest1;

architecture behavior of keybtest1 is

  -- Component Declaration for the Unit Under Test (UUT)
  
  component keyboard
    port(
      reset      : in  std_logic;
      kb_clk     : in  std_logic;
      kb_data    : in  std_logic;
      display    : out std_logic_vector(7 downto 0)
      );
  end component;


  --Inputs
  signal reset   : std_logic := '0';
  signal kb_clk  : std_logic := '0';
  signal kb_data : std_logic := '0';

  --Outputs
  signal display    : std_logic_vector(7 downto 0);

  procedure keyprint (
    constant key     : in  std_logic_vector(7 downto 0);
    signal   kbdata  : out std_logic;
    signal   kbclock : out std_logic) is
  begin  -- keyprint
    -- insert stimulus here 
--    kbclock <= '1';
--    wait for 500 us;
--
--    kbclock <= '0';
--    wait for 65 us;
--    kbclock <= '1';
--    wait for 65 us;

-- start bit
    kbdata  <= '0';
    kbclock <= '0';
    wait for 65 us;
    kbclock <= '1';
    wait for 65 us;

    kbdata  <= key(7);
    kbclock <= '0';
    wait for 65 us;
    kbclock <= '1';
    wait for 65 us;

    kbdata  <= key(6);
    kbclock <= '0';
    wait for 65 us;
    kbclock <= '1';
    wait for 65 us;

    kbdata  <= key(5);
    kbclock <= '0';
    wait for 65 us;
    kbclock <= '1';
    wait for 65 us;

    kbdata  <= key(4);
    kbclock <= '0';
    wait for 65 us;
    kbclock <= '1';
    wait for 65 us;

    kbdata  <= key(3);
    kbclock <= '0';
    wait for 65 us;
    kbclock <= '1';
    wait for 65 us;

    kbdata  <= key(2);
    kbclock <= '0';
    wait for 65 us;
    kbclock <= '1';
    wait for 65 us;

    kbdata  <= key(1);
    kbclock <= '0';
    wait for 65 us;
    kbclock <= '1';
    wait for 65 us;

    kbdata  <= key(0);
    kbclock <= '0';
    wait for 65 us;
    kbclock <= '1';
    wait for 65 us;

-- parity
    kbdata  <= not (key(0) xor key(1) xor key(2) xor key(3) xor key(4) xor key(5) xor key(6) xor key(7));
    kbclock <= '0';
    wait for 65 us;
    kbclock <= '1';
    wait for 65 us;

-- stop bit
    kbdata  <= '1';
    kbclock <= '0';
    wait for 65 us;
    kbclock <= '1';
  end keyprint;

begin

  -- Instantiate the Unit Under Test (UUT)
  uut : keyboard port map (
    reset      => reset,
    kb_clk     => kb_clk,
    kb_data    => kb_data,
    display    => display
    );


  reset_process : process
  begin  -- process reset_process
    wait for 100 ns;
    reset <= '1';
    wait for 100 ns;
    reset <= '0';
    wait;
  end process reset_process;

-- Stimulus process
  stim_proc : process
  begin
    -- hold reset state for 100 ns.
    wait for 1 ms;
    keyprint("10101011", kb_data, kb_clk);
--    wait for 2 ms;
--    keyprint(x"0F", kb_data, kb_clk);
    wait;
  end process;

end;
